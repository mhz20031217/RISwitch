`define IMEM_IMG "/home/pc/Learning/02.IT/5.ICS/ics2023/am-kernels/tests/fpga-tests/build/fpga-tests-riscv32-switch.hex"
`define DMEM_IMG "/home/pc/Learning/02.IT/5.ICS/ics2023/am-kernels/tests/fpga-tests/build/fpga-tests-riscv32-switch_d.hex"
