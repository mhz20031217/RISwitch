`define IMEM_IMG ""
`define DMEM_IMG ""
